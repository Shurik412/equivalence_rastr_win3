JL   `Rastr_for_Win        ���������������info[siga:S,version:I,subversion:I,intcount:I],tabl[namv:S,key:S,desc:S,file:S,tipt:I,fields[name:S,name2:S,tip:I,width:I,prec:I,zag:S,formula:S,afor:I,xrm:I,nameref:S,desc:S,min:D,max:D,mash:D,backr:S,cash:I,redirect:S,exttreex:I,unit:S]]������     #�  �   ,JL
   -D� ������������diff      diff_it      ������� ������������ ����������  !������������ ������.form diff_it tabl col addit vib Xd_a98519 _a98520 _a98521 _a98524 _a185063 ��	�̌���������� ������� ���� � ���������� ������� ���� ��� ��������� ���� �������                                                                                       �?      �?      �?      �?      �?����������耂�퀘����������������è�������������̆р�׆߀����������������info[siga:S,version:I,subversion:I,intcount:I],tabl[namv:S,key:S,desc:S,file:S,tipt:I,fields[name:S,name2:S,tip:I,width:I,prec:I,zag:S,formula:S,afor:I,xrm:I,nameref:S,desc:S,min:D,max:D,mash:D,backr:S,cash:I,redirect:S,exttreex:I,unit:S]],diff[_a98519:I,_a98520:S,_a98521:S,_a98524:S,_a185063:S]��������     P� 5  